* SPICE3 file created from q5b.ext - technology: scmos
.include TSMC_180nm.txt
.param SUPPLY = 1.8
.option scale=0.09u
.global gnd vdd

Vdd vdd gnd 'SUPPLY'

M1000 inv01in a vdd inv00w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1001 inv01in a gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=100 ps=60
M1002 inv02in inv01in vdd inv01w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1003 inv02in inv01in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=100 ps=60
M1004 inv03in inv02in vdd inv02w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1005 inv03in inv02in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=100 ps=60
M1006 inv04in inv03in vdd inv03w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1007 inv04in inv03in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=100 ps=60
M1008 inv05in inv04in vdd inv04w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1009 inv05in inv04in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=100 ps=60
M1010 inv06in inv05in vdd inv05w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1011 inv06in inv05in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=100 ps=60
M1012 inv07in inv06in vdd inv06w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1013 inv07in inv06in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=100 ps=60
M1014 inv08in inv07in vdd inv07w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1015 inv08in inv07in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=100 ps=60
M1016 inv09in inv08in vdd inv08w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1017 inv09in inv08in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=100 ps=60
M1018 inv09out inv09in vdd inv09w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1019 inv09out inv09in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=100 ps=60
M1020 inv011in inv09out vdd inv010w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1021 inv011in inv09out gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=100 ps=60
M1022 inv012in inv011in vdd inv011w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1023 inv012in inv011in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=100 ps=60
M1024 inv013in inv012in vdd inv012w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1025 inv013in inv012in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=100 ps=60
M1026 inv014in inv013in vdd inv013w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1027 inv014in inv013in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=100 ps=60
M1028 inv015in inv014in vdd inv014w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1029 inv015in inv014in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=100 ps=60
M1030 inv10in inv015in vdd inv015w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1031 inv10in inv015in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1032 inv11in inv10in vdd inv10w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1033 inv11in inv10in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1034 inv12in inv11in vdd inv11w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1035 inv12in inv11in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1036 inv13in inv12in vdd inv12w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1037 inv13in inv12in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1038 inv14in inv13in vdd inv13w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1039 inv14in inv13in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1040 inv15in inv14in vdd inv14w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1041 inv15in inv14in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1042 inv16in inv15in vdd inv15w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1043 inv16in inv15in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1044 inv17in inv16in vdd inv16w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1045 inv17in inv16in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1046 inv18in inv17in vdd inv17w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1047 inv18in inv17in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1048 inv19in inv18in vdd inv18w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1049 inv19in inv18in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1050 inv110in inv19in vdd inv19w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1051 inv110in inv19in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1052 inv111in inv110in vdd inv110w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1053 inv111in inv110in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1054 inv112in inv111in vdd inv111w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1055 inv112in inv111in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1056 inv113in inv112in vdd inv112w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1057 inv113in inv112in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1058 inv114in inv113in vdd inv113w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1059 inv114in inv113in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1060 a inv114in vdd inv114w00 CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1061 a inv114in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
C0 inv11in vdd 0.02fF
C1 inv012w00 vdd 0.07fF
C2 vdd inv012in 0.29fF
C3 inv010w00 vdd 0.07fF
C4 inv16in inv15in 0.05fF
C5 inv011in gnd 0.05fF
C6 vdd inv112w00 0.07fF
C7 inv015in gnd 0.13fF
C8 inv08in inv08w00 0.06fF
C9 inv17in inv16in 0.05fF
C10 inv011in vdd 0.02fF
C11 vdd inv113w00 0.07fF
C12 gnd inv113in 0.05fF
C13 vdd inv09w00 0.07fF
C14 inv18in inv17in 0.05fF
C15 vdd inv07in 0.02fF
C16 vdd inv114w00 0.07fF
C17 gnd inv114in 0.05fF
C18 inv12w00 vdd 0.07fF
C19 inv19in inv18in 0.05fF
C20 gnd inv09in 0.05fF
C21 inv04w00 inv04in 0.06fF
C22 inv09out gnd 0.05fF
C23 inv10in vdd 0.02fF
C24 inv110in inv19in 0.05fF
C25 inv011w00 inv012in 0.05fF
C26 gnd inv02in 0.05fF
C27 gnd inv01in 0.13fF
C28 inv111in inv110in 0.05fF
C29 vdd vdd 0.03fF
C30 inv014in vdd 0.29fF
C31 vdd inv06in 0.29fF
C32 vdd inv14in 0.02fF
C33 inv011in inv011w00 0.06fF
C34 vdd inv111w00 0.07fF
C35 inv04w00 vdd 0.07fF
C36 inv11in inv12in 0.05fF
C37 inv10in vdd 0.29fF
C38 vdd inv15in 0.02fF
C39 gnd inv112in 0.05fF
C40 inv00w00 inv01in 0.05fF
C41 vdd inv16in 0.02fF
C42 inv114in inv113in 0.05fF
C43 inv011in inv010w00 0.05fF
C44 gnd inv08in 0.13fF
C45 vdd inv17in 0.02fF
C46 vdd inv07w00 0.07fF
C47 a inv114in 0.05fF
C48 inv12w00 inv13in 0.05fF
C49 inv013w00 vdd 0.07fF
C50 gnd inv014in 0.05fF
C51 vdd inv18in 0.02fF
C52 vdd inv04in 0.02fF
C53 inv10in inv11in 0.05fF
C54 vdd inv19in 0.02fF
C55 a inv01in 0.05fF
C56 vdd inv110in 0.02fF
C57 gnd inv03in 0.05fF
C58 vdd inv01in 0.29fF
C59 vdd vdd 0.03fF
C60 gnd inv015in 0.05fF
C61 vdd inv13w00 0.07fF
C62 inv013in vdd 0.29fF
C63 vdd inv011w00 0.07fF
C64 inv112in inv111in 0.05fF
C65 inv11w00 vdd 0.07fF
C66 inv11in gnd 0.05fF
C67 inv10in inv015w00 0.05fF
C68 vdd vdd 0.03fF
C69 inv113in inv112in 0.05fF
C70 inv12in inv12w00 0.06fF
C71 vdd vdd 0.03fF
C72 vdd inv113in 0.02fF
C73 vdd vdd 0.03fF
C74 inv07in inv07w00 0.06fF
C75 vdd inv114in 0.02fF
C76 inv09out vdd 0.02fF
C77 inv03in vdd 0.29fF
C78 inv05in inv04w00 0.05fF
C79 vdd vdd 0.03fF
C80 gnd inv07in 0.13fF
C81 gnd inv04in 0.05fF
C82 inv10in gnd 0.05fF
C83 inv06in inv05w00 0.05fF
C84 inv03w00 vdd 0.07fF
C85 gnd inv012in 0.05fF
C86 inv015in vdd 0.29fF
C87 vdd vdd 0.03fF
C88 gnd inv13in 0.05fF
C89 vdd vdd 0.03fF
C90 vdd vdd 0.03fF
C91 gnd inv14in 0.13fF
C92 vdd inv111in 0.02fF
C93 inv012w00 inv012in 0.06fF
C94 gnd gnd 0.03fF
C95 inv11w00 inv12in 0.05fF
C96 inv09out inv09in 0.05fF
C97 vdd vdd 0.03fF
C98 inv05in inv04in 0.05fF
C99 inv15w00 inv15in 0.06fF
C100 vdd inv112in 0.02fF
C101 vdd vdd 0.03fF
C102 inv16w00 inv16in 0.06fF
C103 vdd vdd 0.03fF
C104 vdd vdd 0.03fF
C105 inv10in inv10w00 0.06fF
C106 vdd vdd 0.03fF
C107 inv17w00 inv17in 0.06fF
C108 vdd vdd 0.03fF
C109 vdd inv13in 0.29fF
C110 inv03in inv02in 0.05fF
C111 inv05in vdd 0.29fF
C112 inv18w00 inv18in 0.06fF
C113 inv015in inv014in 0.05fF
C114 vdd inv09in 0.02fF
C115 inv19w00 inv19in 0.06fF
C116 gnd gnd 0.03fF
C117 inv09out inv011in 0.05fF
C118 vdd inv04in 0.29fF
C119 inv110w00 inv110in 0.06fF
C120 inv06w00 inv06in 0.06fF
C121 inv013in vdd 0.02fF
C122 inv14w00 inv14in 0.06fF
C123 vdd inv014in 0.02fF
C124 vdd vdd 0.03fF
C125 inv111w00 inv111in 0.06fF
C126 gnd inv15in 0.13fF
C127 vdd vdd 0.03fF
C128 vdd vdd 0.03fF
C129 inv12in vdd 0.02fF
C130 inv03w00 inv03in 0.06fF
C131 gnd inv16in 0.13fF
C132 inv113w00 inv113in 0.06fF
C133 inv10in gnd 0.17fF
C134 gnd inv06in 0.13fF
C135 inv08in vdd 0.29fF
C136 gnd inv17in 0.13fF
C137 inv114w00 inv114in 0.06fF
C138 inv03in inv02w00 0.05fF
C139 gnd inv05in 0.13fF
C140 vdd vdd 0.03fF
C141 gnd inv18in 0.13fF
C142 vdd a 0.52fF IC = 0
C143 inv015in inv014w00 0.05fF
C144 vdd vdd 0.05fF IC = 0
C145 inv09w00 inv09in 0.06fF
C146 gnd inv19in 0.13fF
C147 inv14in inv13in 0.05fF
C148 inv10in inv015in 0.05fF
C149 gnd inv110in 0.13fF
C150 inv06w00 vdd 0.07fF
C151 vdd vdd 0.03fF
C152 inv013in inv012in 0.05fF
C153 vdd inv014w00 0.07fF
C154 gnd inv111in 0.13fF
C155 vdd inv12in 0.29fF
C156 inv112w00 inv112in 0.06fF
C157 vdd inv11in 0.29fF
C158 inv12in inv13in 0.05fF
C159 gnd inv113in 0.13fF
C160 inv08in inv07in 0.05fF
C161 inv03in inv04in 0.05fF
C162 gnd inv114in 0.13fF
C163 inv13in gnd 0.13fF
C164 inv013w00 inv014in 0.05fF
C165 vdd vdd 0.05fF IC = 0
C166 gnd a 0.21fF
C167 gnd inv09in 0.13fF
C168 inv09out gnd 0.13fF
C169 gnd inv01in 0.05fF
C170 inv09out inv010w00 0.06fF
C171 inv06in vdd 0.02fF
C172 gnd inv02in 0.13fF
C173 vdd vdd 0.03fF
C174 vdd inv012in 0.02fF
C175 inv014in inv014w00 0.06fF
C176 inv00w00 a 0.06fF
C177 inv05in vdd 0.02fF
C178 inv01w00 inv01in 0.06fF
C179 inv15in vdd 0.29fF
C180 vdd inv015w00 0.07fF
C181 inv00w00 vdd 0.07fF
C182 gnd inv112in 0.13fF
C183 inv12in gnd 0.05fF
C184 inv02in inv01w00 0.05fF
C185 inv16in vdd 0.29fF
C186 inv011in gnd 0.13fF
C187 gnd inv08in 0.05fF
C188 inv08in inv07w00 0.05fF
C189 vdd inv02in 0.02fF
C190 inv17in vdd 0.29fF
C191 gnd inv014in 0.13fF
C192 inv18in vdd 0.29fF
C193 a vdd 0.02fF
C194 inv19in vdd 0.29fF
C195 inv110in vdd 0.29fF
C196 inv13in inv13w00 0.06fF
C197 inv10w00 vdd 0.07fF
C198 inv111in vdd 0.29fF
C199 gnd inv03in 0.13fF
C200 inv12in gnd 0.13fF
C201 inv01w00 vdd 0.07fF
C202 gnd gnd 0.03fF
C203 inv14in inv13w00 0.05fF
C204 vdd vdd 0.03fF
C205 inv11in gnd 0.13fF
C206 vdd vdd 0.03fF
C207 gnd gnd 0.03fF
C208 inv06w00 inv07in 0.05fF
C209 inv02in inv01in 0.05fF
C210 inv113in vdd 0.29fF
C211 vdd inv02w00 0.07fF
C212 inv114in vdd 0.29fF
C213 gnd inv07in 0.05fF
C214 a vdd 0.29fF
C215 vdd inv09in 0.29fF
C216 gnd inv04in 0.13fF
C217 inv05in inv05w00 0.06fF
C218 inv10w00 inv11in 0.05fF
C219 inv014in inv013in 0.05fF
C220 vdd inv03in 0.02fF
C221 inv01in vdd 0.02fF
C222 inv011in vdd 0.29fF
C223 inv11in inv11w00 0.06fF
C224 vdd vdd 0.03fF
C225 inv06in inv07in 0.05fF
C226 inv02in vdd 0.29fF
C227 gnd gnd 0.03fF
C228 inv16in inv15w00 0.05fF
C229 vdd inv08in 0.02fF
C230 inv02in inv02w00 0.06fF
C231 gnd gnd 0.03fF
C232 inv17in inv16w00 0.05fF
C233 gnd gnd 0.03fF
C234 inv18in inv17w00 0.05fF
C235 inv013w00 inv013in 0.06fF
C236 vdd vdd 0.03fF
C237 inv08in inv09in 0.05fF
C238 gnd gnd 0.03fF
C239 inv19in inv18w00 0.05fF
C240 vdd inv05w00 0.07fF
C241 gnd inv013in 0.13fF
C242 inv015in vdd 0.02fF
C243 gnd gnd 0.02fF
C244 inv110in inv19w00 0.05fF
C245 inv09out vdd 0.29fF
C246 gnd gnd 0.03fF
C247 inv111in inv110w00 0.05fF
C248 inv15in inv14w00 0.05fF
C249 gnd inv14in 0.05fF
C250 vdd vdd 0.03fF
C251 vdd vdd 0.03fF
C252 gnd gnd 0.03fF
C253 inv112in vdd 0.29fF
C254 vdd vdd 0.03fF
C255 inv012w00 inv013in 0.05fF
C256 inv011in inv012in 0.05fF
C257 vdd inv07in 0.29fF
C258 vdd inv15w00 0.07fF
C259 gnd inv15in 0.05fF
C260 gnd gnd 0.03fF
C261 inv113in inv112w00 0.05fF
C262 vdd inv08w00 0.07fF
C263 gnd inv06in 0.05fF
C264 vdd inv16w00 0.07fF
C265 gnd inv16in 0.05fF
C266 gnd gnd 0.03fF
C267 inv114in inv113w00 0.05fF
C268 gnd inv05in 0.05fF
C269 vdd inv17w00 0.07fF
C270 gnd inv17in 0.05fF
C271 gnd inv013in 0.05fF
C272 gnd gnd 0.03fF
C273 a inv114w00 0.05fF
C274 vdd inv13in 0.02fF
C275 inv08w00 inv09in 0.05fF
C276 vdd inv18w00 0.07fF
C277 gnd inv18in 0.05fF
C278 inv015in inv015w00 0.06fF
C279 vdd inv19w00 0.07fF
C280 gnd inv19in 0.05fF
C281 inv09out inv09w00 0.05fF
C282 gnd gnd 0.03fF
C283 vdd inv14in 0.29fF
C284 vdd inv110w00 0.07fF
C285 gnd inv110in 0.05fF
C286 gnd inv012in 0.13fF
C287 vdd vdd 0.03fF
C288 inv05in inv06in 0.05fF
C289 inv03w00 inv04in 0.05fF
C290 vdd inv14w00 0.07fF
C291 inv15in inv14in 0.05fF
C292 inv112in inv111w00 0.05fF
C293 gnd inv111in 0.05fF
C294 vdd Gnd 0.55fF 
C295 gnd Gnd 0.23fF
C296 a Gnd 0.41fF
C297 vdd Gnd 0.05fF
C298 inv114w00 Gnd 0.89fF
C299 gnd Gnd 0.23fF
C300 inv114in Gnd 0.22fF
C301 vdd Gnd 0.05fF
C302 inv113w00 Gnd 0.89fF
C303 gnd Gnd 0.23fF
C304 inv113in Gnd 0.22fF
C305 vdd Gnd 0.05fF
C306 inv112w00 Gnd 0.89fF
C307 gnd Gnd 0.23fF
C308 inv112in Gnd 0.22fF
C309 vdd Gnd 0.05fF
C310 inv111w00 Gnd 0.89fF
C311 gnd Gnd 0.23fF
C312 inv111in Gnd 0.22fF
C313 vdd Gnd 0.05fF
C314 inv110w00 Gnd 0.89fF
C315 gnd Gnd 0.23fF
C316 inv110in Gnd 0.22fF
C317 vdd Gnd 0.05fF
C318 inv19w00 Gnd 0.89fF
C319 gnd Gnd 0.23fF
C320 inv19in Gnd 0.22fF
C321 vdd Gnd 0.05fF
C322 inv18w00 Gnd 0.89fF
C323 gnd Gnd 0.23fF
C324 inv18in Gnd 0.22fF
C325 vdd Gnd 0.05fF
C326 inv17w00 Gnd 0.89fF
C327 gnd Gnd 0.23fF
C328 inv17in Gnd 0.22fF
C329 vdd Gnd 0.05fF
C330 inv16w00 Gnd 0.89fF
C331 gnd Gnd 0.23fF
C332 inv16in Gnd 0.22fF
C333 vdd Gnd 0.05fF
C334 inv15w00 Gnd 0.89fF
C335 gnd Gnd 0.23fF
C336 inv15in Gnd 0.22fF
C337 vdd Gnd 0.05fF
C338 inv14w00 Gnd 0.89fF
C339 gnd Gnd 0.23fF
C340 inv14in Gnd 0.22fF
C341 vdd Gnd 0.05fF
C342 inv13w00 Gnd 0.89fF
C343 gnd Gnd 0.23fF
C344 inv13in Gnd 0.22fF
C345 vdd Gnd 0.05fF
C346 inv12w00 Gnd 0.89fF
C347 gnd Gnd 0.23fF
C348 inv12in Gnd 0.22fF
C349 vdd Gnd 0.05fF
C350 inv11w00 Gnd 0.89fF
C351 gnd Gnd 0.23fF
C352 inv11in Gnd 0.22fF
C353 vdd Gnd 0.05fF
C354 inv10in Gnd 0.49fF
C355 inv10w00 Gnd 0.89fF
C356 gnd Gnd 0.12fF
C357 vdd Gnd 0.05fF
C358 inv015in Gnd 0.22fF
C359 inv015w00 Gnd 0.89fF
C360 vdd Gnd 0.05fF
C361 inv014in Gnd 0.22fF
C362 inv014w00 Gnd 0.89fF
C363 vdd Gnd 0.05fF
C364 inv013in Gnd 0.22fF
C365 inv013w00 Gnd 0.89fF
C366 vdd Gnd 0.05fF
C367 inv012in Gnd 0.22fF
C368 inv012w00 Gnd 0.89fF
C369 vdd Gnd 0.05fF
C370 inv011in Gnd 0.22fF
C371 inv011w00 Gnd 0.89fF
C372 vdd Gnd 0.05fF
C373 inv09out Gnd 0.22fF
C374 inv010w00 Gnd 0.89fF
C375 vdd Gnd 0.05fF
C376 inv09in Gnd 0.22fF
C377 inv09w00 Gnd 0.89fF
C378 vdd Gnd 0.05fF
C379 inv08in Gnd 0.22fF
C380 inv08w00 Gnd 0.89fF
C381 vdd Gnd 0.05fF
C382 inv07in Gnd 0.22fF
C383 inv07w00 Gnd 0.89fF
C384 vdd Gnd 0.05fF
C385 inv06in Gnd 0.22fF
C386 inv06w00 Gnd 0.89fF
C387 vdd Gnd 0.05fF
C388 inv05in Gnd 0.22fF
C389 inv05w00 Gnd 0.89fF
C390 vdd Gnd 0.05fF
C391 inv04in Gnd 0.22fF
C392 inv04w00 Gnd 0.89fF
C393 vdd Gnd 0.05fF
C394 inv03in Gnd 0.22fF
C395 inv03w00 Gnd 0.89fF
C396 vdd Gnd 0.05fF
C397 inv02in Gnd 0.22fF
C398 inv02w00 Gnd 0.89fF
C399 vdd Gnd 0.05fF
C400 inv01in Gnd 0.22fF
C401 inv01w00 Gnd 0.89fF
C402 vdd Gnd 0.05fF
C403 inv00w00 Gnd 0.89fF
.ic v(a) 1.8
.tran 10p 10n
.measure tran tperiod
+ TRIG v(a) VAL='SUPPLY/2' RISE=1
+ TARG v(a) VAL='SUPPLY/2' RISE=2
.control
set hcopypscolor = 1 *White background for saving plots
set color0=white 
set color1=black 

run
set curplottitle= "siva-2019102038-5-b"
plot v(a)
.endc
.end
